class Instruction;
   rand bit [15:0] Instr;
endclass; // Instruction
