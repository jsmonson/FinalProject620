package EnvironmentPkg;

`include "Instruction.sv"
`include "ScoreBoard.sv"
   
endpackage