class Scoreboard;

endclass // Scoreboard
